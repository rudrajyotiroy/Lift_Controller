// This file should be compile top spec (temporarily)

`include "lift_controller_if.sv"
`include "request_handler.v"
`include "door_controller.v"
`include "main_alu_block.v"
`include "lift_controller_wrapper.v"
`include "lift_movement_emulator.sv"
`include "tb_top.sv"