`ifndef LIFT_CONTROLLER_DEFINES
`define LIFT_CONTROLLER_DEFINES

`define MAX_REQUESTS 20
`define NUM_FLOORS 12
`define DRAIN_TIME 50000

`endif