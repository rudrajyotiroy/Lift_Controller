`ifndef LIFT_CONTROLLER_DEFINES
`define LIFT_CONTROLLER_DEFINES

`define MAX_REQUESTS 100
`define NUM_FLOORS 24
`define DRAIN_TIME 500000

`define MONO_LIFT
`define DEBUG_INTERFACE

`endif